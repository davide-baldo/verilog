`ifndef _H_CLOCK_
`define _H_CLOCK_

interface Clock;
  logic stop_clock;
  wire signal;
endinterface

`endif /* _H_CLOCK_ */