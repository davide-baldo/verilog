`ifndef _H_CONF_
`define _H_CONF_

`define ARCH_SIZE 64

`define ARCH_SIZE_1 63

/* verilator lint_off CASEINCOMPLETE */
/* verilator lint_off WIDTH */

`endif /* _H_CONF_ */