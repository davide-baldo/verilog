`ifndef _H_CONF_
`define _H_CONF_

`define ARCH_SIZE 64

`define ARCH_SIZE_1 63

`endif /* _H_CONF_ */